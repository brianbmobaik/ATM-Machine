`timescale 1ns / 1ps

module BtnUpDown (
    input wire rst,
    input wire [1:0] UpDown,
    output reg [3:0] data
    );
endmodule