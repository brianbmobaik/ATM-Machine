`timescale 1ns/1ps

module TestModule (
    input clk, rst,
    input [4:0] btn,
    input 
    );

    
endmodule