`timescale 1ns / 1ps

module BtnLeftRight ();
endmodule